module main(a,b);
input a;output b;output c; output d;
assign b=a;
assign c=a;
assign d=a;
endmodule
module main(a,b);
input a;output b;output c;
assign b=a;
assign c=a;
endmodule
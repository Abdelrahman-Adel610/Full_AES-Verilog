`include "InvShiftRows.v"
`include "InvSubBytes.v"
`include "Inv_MixColumns.v"
`include "AddRoundKey.v"
module DecryptionRound(
    input wire [127:0] instate,
    input wire [127:0] roundKey,	
    output wire [127:0] outstate
);
wire [127:0] InvSubBytes_outstate;
wire [127:0] InvShiftRows_outstate;
wire [127:0] Inv_MixColumns_outstate;
wire [127:0] AddRoundKey_outstate;
assign instate=128'h193de3bea0f4e22b9ac68d2aeaf84808;
assign roundKey=128'hac7766f319fadc2128d12941575c006a;
InvSubBytes  op1 (instate,InvSubBytes_outstate);
InvShiftRows  op2 (InvSubBytes_outstate,InvShiftRows_outstate);
AddRoundKey op3 (InvShiftRows_outstate,AddRoundKey_outstate, );
Inv_MixColumns  op4 (AddRoundKey_outstate,Inv_MixColumns_outstate);
assign outstate=Inv_MixColumns_outstate;
endmodule
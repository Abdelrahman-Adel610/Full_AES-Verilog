`include "EncryptionRound.v"
`include "DecryptionRound.v"


module main(
    input wire [127:0] instate,	
    output wire [127:0] outstate
);

endmodule
 //Testbench
module Test_ShiftRows();

reg [127:0] in;
wire [127:0] out;

initial begin
    in = 128'h3243f6a8885a308d313198a2e0370734;
end

ShiftRows test(in, out);

endmodule
//Testbench:
module Test_InvShiftRows();

reg [127:0] in;
wire [127:0] out;

initial begin
    in = 128'h325a9834883107a83137f68de04330a2;
end

InvShiftRows test(in, out);

endmodule
`include "EncryptionRound.v"
`include "InvShiftRows.v"
`include "InvSubBytes.v"
`include "Inv_MixColumns.v"

module main(
    input wire [127:0] instate,	
    output wire [127:0] outstate
);

endmodule
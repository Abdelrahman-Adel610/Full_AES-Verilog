`include "ShiftRows.v"
`include "SubBytes.v"
`include "InvShiftRows.v"
`include "InvSubBytes.v"
module main;

endmodule
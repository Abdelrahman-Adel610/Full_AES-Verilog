module main(a,b);
input a;output b;output d;
assign b=a;
endmodule
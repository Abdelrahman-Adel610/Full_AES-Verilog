`include "InvShiftRows.v"
`include "InvSubBytes.v"
`include "Inv_MixColumns.v"
`include "AddRoundKey.v"
`include "DecryptionRound.v"
`include "KeyExpansion.v"
module AES_Decryption(input [127:0] in , output [127:0] out , input [127:0] Key, input clk);
wire [1407:0] state;
wire [1407:0] full_key;
wire [127:0] InvSubBytes_out;
wire [127:0] InvShiftRows_out;
reg[3:0] i;
initial i=0;
DecryptionRound dr (state[(i*(-128)+1407)-:128] , full_key [(i*(-128)+1407)-:128] ,state[(i*(-128)+1279)-:128]);   	
always @(posedge clk)
begin
   if (i<10)
    begin   

        i=i+1;
   end
end


KeyExpansion kr(Key , full_key);  
 AddRoundKey preak (in , InvSubBytes_out , full_key[1407-:128]);
 InvShiftRows preIsh (InvSubBytes_out , InvShiftRows_out);
 InvSubBytes preIsu (InvShiftRows_out , state[1279-:128]);
 /*
genvar i;
generate
    for (i = 1 ; i < 10 ; i = i + 1 ) begin : decryp
      	DecryptionRound dr (state[(i*(-128)+1407)-:128] , full_key [(i*(-128)+1407)-:128] ,state[(i*(-128)+1279)-:128] , clk); // in , key , out
      	// $monitor(?Time=%0d state[(i*(-128)+1535)-:128]=%b full_key [(i*(-128)+1407)-:128]=%b state[(i*(-128)+1407)-:128]=%b?, $time,state[(i*(-128)+1535)-:128],full_key [(i*(-128)+1407)-:128],state[(i*(-128)+1407)-:128]);
    end
endgenerate*/
  AddRoundKey ak (state[127:0] ,out ,full_key[127:0]);


/*
always@( posedge clk) begin
 out <= state[127:0];
end*/
endmodule